// Copyright Supranational LLC
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

    MINROOT_VDF_CONTROL = csr_addr_t'('h200000),//csr-pkg-include
    MINROOT_VDF_CMD_JOB_ID = csr_addr_t'('h201000),//csr-pkg-include
    MINROOT_VDF_CMD_ITER_COUNT_0 = csr_addr_t'('h201004),//csr-pkg-include
    MINROOT_VDF_CMD_ITER_COUNT_1 = csr_addr_t'('h201008),//csr-pkg-include
    MINROOT_VDF_CMD_START_ITER_0 = csr_addr_t'('h20100c),//csr-pkg-include
    MINROOT_VDF_CMD_START_ITER_1 = csr_addr_t'('h201010),//csr-pkg-include
    MINROOT_VDF_CMD_X_0 = csr_addr_t'('h201014),//csr-pkg-include
    MINROOT_VDF_CMD_X_1 = csr_addr_t'('h201018),//csr-pkg-include
    MINROOT_VDF_CMD_X_2 = csr_addr_t'('h20101c),//csr-pkg-include
    MINROOT_VDF_CMD_X_3 = csr_addr_t'('h201020),//csr-pkg-include
    MINROOT_VDF_CMD_X_4 = csr_addr_t'('h201024),//csr-pkg-include
    MINROOT_VDF_CMD_X_5 = csr_addr_t'('h201028),//csr-pkg-include
    MINROOT_VDF_CMD_X_6 = csr_addr_t'('h20102c),//csr-pkg-include
    MINROOT_VDF_CMD_X_7 = csr_addr_t'('h201030),//csr-pkg-include
    MINROOT_VDF_CMD_X_8 = csr_addr_t'('h201034),//csr-pkg-include
    MINROOT_VDF_CMD_X_9 = csr_addr_t'('h201038),//csr-pkg-include
    MINROOT_VDF_CMD_Y_0 = csr_addr_t'('h20103c),//csr-pkg-include
    MINROOT_VDF_CMD_Y_1 = csr_addr_t'('h201040),//csr-pkg-include
    MINROOT_VDF_CMD_Y_2 = csr_addr_t'('h201044),//csr-pkg-include
    MINROOT_VDF_CMD_Y_3 = csr_addr_t'('h201048),//csr-pkg-include
    MINROOT_VDF_CMD_Y_4 = csr_addr_t'('h20104c),//csr-pkg-include
    MINROOT_VDF_CMD_Y_5 = csr_addr_t'('h201050),//csr-pkg-include
    MINROOT_VDF_CMD_Y_6 = csr_addr_t'('h201054),//csr-pkg-include
    MINROOT_VDF_CMD_Y_7 = csr_addr_t'('h201058),//csr-pkg-include
    MINROOT_VDF_CMD_Y_8 = csr_addr_t'('h20105c),//csr-pkg-include
    MINROOT_VDF_CMD_Y_9 = csr_addr_t'('h201060),//csr-pkg-include
    MINROOT_VDF_CMD_START = csr_addr_t'('h201064),//csr-pkg-include
    MINROOT_VDF_STATUS_JOB_ID = csr_addr_t'('h202000),//csr-pkg-include
    MINROOT_VDF_STATUS_ITER_0 = csr_addr_t'('h202004),//csr-pkg-include
    MINROOT_VDF_STATUS_ITER_1 = csr_addr_t'('h202008),//csr-pkg-include
    MINROOT_VDF_STATUS_X_0 = csr_addr_t'('h20200c),//csr-pkg-include
    MINROOT_VDF_STATUS_X_1 = csr_addr_t'('h202010),//csr-pkg-include
    MINROOT_VDF_STATUS_X_2 = csr_addr_t'('h202014),//csr-pkg-include
    MINROOT_VDF_STATUS_X_3 = csr_addr_t'('h202018),//csr-pkg-include
    MINROOT_VDF_STATUS_X_4 = csr_addr_t'('h20201c),//csr-pkg-include
    MINROOT_VDF_STATUS_X_5 = csr_addr_t'('h202020),//csr-pkg-include
    MINROOT_VDF_STATUS_X_6 = csr_addr_t'('h202024),//csr-pkg-include
    MINROOT_VDF_STATUS_X_7 = csr_addr_t'('h202028),//csr-pkg-include
    MINROOT_VDF_STATUS_X_8 = csr_addr_t'('h20202c),//csr-pkg-include
    MINROOT_VDF_STATUS_X_9 = csr_addr_t'('h202030),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_0 = csr_addr_t'('h202034),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_1 = csr_addr_t'('h202038),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_2 = csr_addr_t'('h20203c),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_3 = csr_addr_t'('h202040),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_4 = csr_addr_t'('h202044),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_5 = csr_addr_t'('h202048),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_6 = csr_addr_t'('h20204c),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_7 = csr_addr_t'('h202050),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_8 = csr_addr_t'('h202054),//csr-pkg-include
    MINROOT_VDF_STATUS_Y_9 = csr_addr_t'('h202058),//csr-pkg-include
    MINROOT_VDF_STATUS_END = csr_addr_t'('h20205c),//csr-pkg-include
    MINROOT_VDF_RW = csr_addr_t'('h20fff8),//csr-pkg-include
    MINROOT_VDF_END_OF_RANGE = csr_addr_t'('h20fffc)//csr-pkg-include
